// windowBuffer.v
// Adaptive Median Filter
// Windows Buffer module
// AUTHOR : Reza Bahrami
// Email : r.bahrami.work@outlook.com

// MIT License
// 
// Copyright (c) 2021 Reza Bahrami
// 
// Permission is hereby granted, free of charge, to any person obtaining a copy
// of this software and associated documentation files (the "Software"), to deal
// in the Software without restriction, including without limitation the rights
// to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
// copies of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:
// 
// The above copyright notice and this permission notice shall be included in all
// copies or substantial portions of the Software.
// 
// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
// IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
// FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
// AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
// LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
// OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
// SOFTWARE.

`default_nettype none

module windowBuffer (out, wCenter, in, windowF);
	// Parameters
	parameter WINDOW_BITS = 200, DATA_WIDTH = 8, CENTER = 12;
	// Outputs
	output reg [WINDOW_BITS - 1 : 0] 		out;
	output reg [DATA_WIDTH - 1 : 0]	wCenter;
	// Inputs
	input wire [WINDOW_BITS - 1 : 0] in;
	input wire windowF;

	// Behavioral Description of module
	always @(posedge windowF) begin
		out = in;
		wCenter = in[(DATA_WIDTH * CENTER + (DATA_WIDTH - 1)) : (DATA_WIDTH * CENTER)];
	end
endmodule