// sram.v
// Adaptive Median Filter
// SRAM Module
// AUTHOR : Reza Bahrami
// Email : r.bahrami.work@outlook.com

// MIT License
// 
// Copyright (c) 2021 Reza Bahrami
// 
// Permission is hereby granted, free of charge, to any person obtaining a copy
// of this software and associated documentation files (the "Software"), to deal
// in the Software without restriction, including without limitation the rights
// to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
// copies of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:
// 
// The above copyright notice and this permission notice shall be included in all
// copies or substantial portions of the Software.
// 
// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
// IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
// FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
// AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
// LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
// OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
// SOFTWARE.

`default_nettype none

module sram (dataOut, dataIn, addr, wr, clk, rst);
	// Parameters
	parameter ADDR_WIDTH = 8, DATA_WIDTH = 8, DEPTH = 256;
	
	// I/Os
	output reg [DATA_WIDTH - 1 : 0] dataOut;
	input wire [DATA_WIDTH - 1 : 0] dataIn;
	input wire [ADDR_WIDTH - 1 : 0] addr;
	input wire wr, clk, rst;

	// Internal Registers
	reg [DATA_WIDTH - 1 : 0] mem [DEPTH - 1 : 0];

	// Module Behavioral Description
	always @(negedge clk)
		if(wr) mem[addr] <= dataIn;
		else dataOut <= mem[addr];

	integer index;
	always @(posedge rst)
		for (index = 0; index < DEPTH; index = index + 1)
			mem[index] <= 0;
endmodule